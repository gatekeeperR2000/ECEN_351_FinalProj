*******************************************************************************
* CDL netlist
*
* Library : Final
* Top Cell Name: Register_File
* View Name: extracted
* Netlist created: 03.Apr.2023 13:05:14
*******************************************************************************

*.SCALE METER
.GLOBAL vdd
.GLOBAL vss

*******************************************************************************
* Library Name: Final
* Cell Name:    Register_File
* View Name:    extracted
*******************************************************************************

.SUBCKT Register_File Addr0 Addr1 Addr2
*.PININFO Addr0:B Addr1:B Addr2:B

MM248 n120 n14 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.35e-06 $Y=7.35e-05
MM0 n93 Addr0 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-3.885e-05 $Y=0.0001821
MM389 n4 Addr0 n147 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001194 $Y=7.35e-05
MM106 n140 n35 n151 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.965e-05 $Y=3.3e-06
MM281 n4 n10 n138 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.505e-05 $Y=6.33e-05
MM128 n165 n76 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.435e-05 $Y=5.01e-05
MM212 n4 n96 n71 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.965e-05 $Y=0.0001671
MM340 n58 n139 n90 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.945e-05 $Y=0.0001671
MM198 n27 n147 n172 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001593 $Y=8.85e-05
MM152 n3 n173 n61 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.905e-05 $Y=5.01e-05
MM236 n169 n71 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.65e-06 $Y=0.0001671
MM291 n140 n175 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.015e-05 $Y=1.65e-05
MM311 n74 n99 n5 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.965e-05 $Y=0.0001101
MM301 n4 n15 n131 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.455e-05 $Y=0.0001569
MM35 n142 n169 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.35e-06 $Y=0.0001821
MM257 n4 n155 n114 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.245e-05 $Y=6.33e-05
MM276 n23 n144 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.505e-05 $Y=0.0001671
MM210 n96 Addr1 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-3.885e-05 $Y=0.0001569
MM338 n28 n45 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.435e-05 $Y=2.67e-05
MM75 n162 n23 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.015e-05 $Y=0.0001821
MM34 n179 n19 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-7.65e-06 $Y=3.3e-06
MM204 n3 n101 n100 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001884 $Y=9.69e-05
MM266 n123 n57 n17 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.755e-05 $Y=2.67e-05
MM61 n127 n29 n51 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.995e-05 $Y=0.0001353
MM219 n19 Addr2 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.965e-05 $Y=1.65e-05
MM4 n3 n111 n91 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.965e-05 $Y=0.0001437
MM356 n4 n58 n109 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.905e-05 $Y=0.0001671
MM30 n157 n33 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-7.65e-06 $Y=9.69e-05
MM357 n115 n153 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.905e-05 $Y=0.0001569
MM290 n4 n36 n41 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.015e-05 $Y=2.67e-05
MM268 n154 n37 n144 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.995e-05 $Y=0.0001671
MM174 n3 n88 n128 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.435e-05 $Y=9.69e-05
MM76 n55 n121 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.015e-05 $Y=0.0001437
MM310 n26 n59 n38 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.965e-05 $Y=0.0001203
MM7 n156 Addr1 n3 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.965e-05 $Y=8.49e-05
MM252 n37 n142 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.245e-05 $Y=0.0001671
MM207 n105 n177 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000201 $Y=9.69e-05
MM196 n50 n161 n172 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001569 $Y=8.85e-05
MM352 n18 n8 n92 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.185e-05 $Y=7.35e-05
MM396 n166 n47 n52 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001419 $Y=0.0001101
MM18 n104 n93 n182 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.725e-05 $Y=3.3e-06
MM374 n69 n22 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.925e-05 $Y=0.0001203
MM282 n4 n123 n36 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.505e-05 $Y=2.67e-05
MM250 n57 n183 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.35e-06 $Y=2.67e-05
MM130 n3 n7 n20 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.435e-05 $Y=3.3e-06
MM217 n75 Addr2 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.965e-05 $Y=6.33e-05
MM317 n42 n15 n86 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.205e-05 $Y=0.0001569
MM28 n3 n16 n129 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-7.65e-06 $Y=0.0001437
MM12 n79 Addr0 n91 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.725e-05 $Y=0.0001437
MM235 n19 n96 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.485e-05 $Y=1.65e-05
MM170 n3 n167 n63 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.925e-05 $Y=3.3e-06
MM175 n27 n130 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.435e-05 $Y=8.85e-05
MM39 n3 n14 n120 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.35e-06 $Y=8.85e-05
MM331 n7 n151 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.925e-05 $Y=1.65e-05
MM60 n64 n53 n52 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.995e-05 $Y=0.0001437
MM136 n76 n135 n173 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.945e-05 $Y=5.01e-05
MM133 n159 n59 n66 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.945e-05 $Y=0.0001353
MM297 n30 n21 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.945e-05 $Y=6.33e-05
MM305 n4 n30 n135 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.455e-05 $Y=6.33e-05
MM300 n4 n139 n46 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.455e-05 $Y=0.0001671
MM80 n132 n138 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.015e-05 $Y=5.01e-05
MM172 n52 n158 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.435e-05 $Y=0.0001437
MM167 n130 n12 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.925e-05 $Y=8.85e-05
MM336 n110 n125 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.435e-05 $Y=7.35e-05
MM193 n24 n178 n65 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001518 $Y=9.69e-05
MM64 n10 n155 n50 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.995e-05 $Y=5.01e-05
MM372 n149 n109 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.925e-05 $Y=0.0001671
MM140 n153 n15 n95 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.185e-05 $Y=0.0001437
MM354 n122 n85 n60 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.185e-05 $Y=2.67e-05
MM17 n9 Addr0 n108 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.725e-05 $Y=3.81e-05
MM178 n78 n63 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.435e-05 $Y=3.3e-06
MM124 n3 n72 n86 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.435e-05 $Y=0.0001437
MM90 n3 n21 n35 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.945e-05 $Y=3.3e-06
MM165 n69 n22 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.925e-05 $Y=0.0001353
MM187 n166 n67 n52 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001419 $Y=9.69e-05
MM367 n136 n39 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.415e-05 $Y=0.0001101
MM154 n167 n77 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.905e-05 $Y=3.3e-06
MM320 n73 n87 n110 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.205e-05 $Y=7.35e-05
MM27 n169 n71 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-7.65e-06 $Y=0.0001821
MM67 n23 n144 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.505e-05 $Y=0.0001821
MM205 n107 n100 n177 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001935 $Y=9.69e-05
MM203 n3 Addr2 n101 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001833 $Y=9.69e-05
MM20 n16 n96 n79 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.485e-05 $Y=0.0001437
MM233 n75 Addr1 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.485e-05 $Y=6.33e-05
MM220 n4 n93 n71 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.725e-05 $Y=0.0001671
MM360 n12 n92 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.905e-05 $Y=7.35e-05
MM415 n54 n100 n177 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001959 $Y=0.0001101
MM82 n140 n175 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.015e-05 $Y=3.3e-06
MM164 n158 n115 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.925e-05 $Y=0.0001437
MM359 n4 n164 n39 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.905e-05 $Y=0.0001101
MM59 n154 n142 n144 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.995e-05 $Y=0.0001821
MM386 n4 n124 n25 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.435e-05 $Y=2.67e-05
MM31 n14 n116 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-7.65e-06 $Y=8.85e-05
MM72 n3 n10 n138 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.505e-05 $Y=5.01e-05
MM221 n4 Addr0 n16 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.725e-05 $Y=0.0001569
MM369 n44 n61 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.415e-05 $Y=6.33e-05
MM150 n39 n164 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.905e-05 $Y=9.69e-05
MM273 n10 n114 n50 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.995e-05 $Y=6.33e-05
MM73 n36 n123 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.505e-05 $Y=4.17e-05
MM238 n49 n103 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.65e-06 $Y=0.0001203
MM365 n4 n115 n95 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.415e-05 $Y=0.0001569
MM127 n3 n125 n110 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.435e-05 $Y=8.85e-05
MM46 n3 n137 n150 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.245e-05 $Y=9.69e-05
MM48 n3 n155 n114 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.245e-05 $Y=5.01e-05
MM173 n3 n69 n51 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.435e-05 $Y=0.0001353
MM370 n122 n6 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.415e-05 $Y=2.67e-05
MM186 n3 n62 n32 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001347 $Y=8.85e-05
MM309 n42 n131 n55 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.965e-05 $Y=0.0001569
MM308 n152 n46 n162 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.965e-05 $Y=0.0001671
MM211 n4 Addr2 n111 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-3.885e-05 $Y=0.0001203
MM137 n45 n85 n60 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.945e-05 $Y=4.17e-05
MM58 n89 n145 n17 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.755e-05 $Y=3.3e-06
MM255 n150 n137 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.245e-05 $Y=0.0001101
MM295 n84 n21 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.945e-05 $Y=0.0001101
MM66 n78 n81 n89 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.995e-05 $Y=3.3e-06
MM397 n25 n161 n82 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001419 $Y=7.35e-05
MM316 n152 n139 n126 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.205e-05 $Y=0.0001671
MM199 n3 n65 n11 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001665 $Y=9.69e-05
MM227 n4 n93 n19 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.725e-05 $Y=1.65e-05
MM131 n58 n46 n90 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.945e-05 $Y=0.0001821
MM32 n171 n75 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-7.65e-06 $Y=5.01e-05
MM225 n75 n93 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.725e-05 $Y=6.33e-05
MM385 n4 n68 n50 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.435e-05 $Y=6.33e-05
MM280 n4 n56 n133 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.505e-05 $Y=7.35e-05
MM25 n43 Addr2 n108 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.485e-05 $Y=3.81e-05
MM344 n92 n87 n125 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.945e-05 $Y=7.35e-05
MM303 n4 n84 n99 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.455e-05 $Y=0.0001101
MM269 n64 n119 n52 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.995e-05 $Y=0.0001569
MM339 n20 n7 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.435e-05 $Y=1.65e-05
MM394 n141 n178 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001347 $Y=0.0001101
MM353 n173 n135 n44 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.185e-05 $Y=6.33e-05
MM246 n29 n49 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.35e-06 $Y=0.0001203
MM99 n152 n139 n162 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.965e-05 $Y=0.0001821
MM403 n94 n32 n172 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001518 $Y=7.35e-05
MM299 n4 n21 n35 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.945e-05 $Y=1.65e-05
MM141 n66 n97 n112 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.185e-05 $Y=0.0001353
MM177 n25 n124 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.435e-05 $Y=4.17e-05
MM53 n127 n40 n17 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.755e-05 $Y=0.0001353
MM241 n4 n75 n171 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.65e-06 $Y=6.33e-05
MM322 n28 n83 n48 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.205e-05 $Y=2.67e-05
MM215 n4 n111 n33 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.965e-05 $Y=0.0001101
MM329 n4 n106 n76 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.925e-05 $Y=6.33e-05
MM78 n5 n98 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.015e-05 $Y=9.69e-05
MM8 n148 Addr2 n3 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.965e-05 $Y=5.01e-05
MM287 n4 n98 n5 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.015e-05 $Y=0.0001101
MM162 n143 n167 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.415e-05 $Y=3.3e-06
MM190 n78 n161 n82 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001443 $Y=8.85e-05
MM10 n3 Addr2 n182 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.965e-05 $Y=3.3e-06
MM13 n134 n93 n163 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.725e-05 $Y=0.0001317
MM195 n24 n47 n51 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001569 $Y=9.69e-05
MM201 n3 n11 n54 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001716 $Y=9.69e-05
MM229 n16 n96 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.485e-05 $Y=0.0001569
MM230 n103 n111 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.485e-05 $Y=0.0001203
MM231 n4 Addr1 n33 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.485e-05 $Y=0.0001101
MM362 n6 n60 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.905e-05 $Y=2.67e-05
MM96 n3 n30 n135 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.455e-05 $Y=5.01e-05
MM116 n3 n42 n72 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.925e-05 $Y=0.0001437
MM145 n122 n83 n60 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.185e-05 $Y=4.17e-05
MM315 n140 n80 n151 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.965e-05 $Y=1.65e-05
MM77 n38 n70 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.015e-05 $Y=0.0001353
MM143 n18 n87 n92 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.185e-05 $Y=8.85e-05
MM91 n3 n139 n46 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.455e-05 $Y=0.0001821
MM412 n4 Addr2 n101 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001833 $Y=0.0001101
MM355 n143 n80 n77 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.185e-05 $Y=1.65e-05
MM313 n106 n135 n132 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.965e-05 $Y=6.33e-05
MM179 n3 Addr0 n67 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001194 $Y=9.69e-05
MM63 n56 n120 n27 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.995e-05 $Y=8.85e-05
MM33 n183 n43 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-7.65e-06 $Y=4.17e-05
MM92 n3 n15 n131 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.455e-05 $Y=0.0001437
MM44 n119 n53 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.245e-05 $Y=0.0001437
MM399 n78 n147 n82 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001443 $Y=7.35e-05
MM87 n87 n21 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.945e-05 $Y=8.85e-05
MM181 n3 Addr1 n178 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001245 $Y=9.69e-05
MM166 n3 n39 n88 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.925e-05 $Y=9.69e-05
MM390 n178 Addr1 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001245 $Y=0.0001101
MM325 n4 n42 n72 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.925e-05 $Y=0.0001569
MM5 n134 Addr1 n3 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.965e-05 $Y=0.0001317
MM109 n26 n59 n31 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.205e-05 $Y=0.0001353
MM261 n64 n53 n17 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.755e-05 $Y=0.0001569
MM226 n4 Addr0 n43 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.725e-05 $Y=2.67e-05
MM21 n103 n111 n163 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.485e-05 $Y=0.0001317
MM119 n3 n73 n125 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.925e-05 $Y=8.85e-05
MM407 n27 n161 n172 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001593 $Y=7.35e-05
MM142 n136 n84 n164 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.185e-05 $Y=9.69e-05
MM94 n3 n84 n99 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.455e-05 $Y=9.69e-05
MM364 n4 n109 n34 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.415e-05 $Y=0.0001671
MM112 n106 n135 n165 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.205e-05 $Y=5.01e-05
MM19 n71 n111 n160 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.485e-05 $Y=0.0001785
MM148 n3 n153 n115 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.905e-05 $Y=0.0001437
MM306 n4 n83 n85 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.455e-05 $Y=2.67e-05
MM240 n14 n116 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.65e-06 $Y=7.35e-05
MM89 n83 n21 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.945e-05 $Y=4.17e-05
MM70 n3 n146 n98 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.505e-05 $Y=9.69e-05
MM333 n86 n72 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.435e-05 $Y=0.0001569
MM68 n3 n64 n121 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.505e-05 $Y=0.0001437
MM382 n51 n69 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.435e-05 $Y=0.0001203
MM327 n4 n74 n118 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.925e-05 $Y=0.0001101
MM289 n132 n138 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.015e-05 $Y=6.33e-05
MM50 n145 n81 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.245e-05 $Y=3.3e-06
MM319 n74 n84 n13 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.205e-05 $Y=0.0001101
MM153 n6 n60 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.905e-05 $Y=4.17e-05
MM406 n24 n47 n128 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001593 $Y=0.0001101
MM249 n4 n171 n155 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.35e-06 $Y=6.33e-05
MM85 n97 n21 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.945e-05 $Y=0.0001353
MM191 n166 n141 n65 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001494 $Y=9.69e-05
MM368 n4 n12 n18 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.415e-05 $Y=7.35e-05
MM383 n128 n88 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.435e-05 $Y=0.0001101
MM377 n68 n61 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.925e-05 $Y=6.33e-05
MM243 n179 n19 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.65e-06 $Y=1.65e-05
MM139 n34 n139 n58 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.185e-05 $Y=0.0001821
MM228 n71 n111 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.485e-05 $Y=0.0001671
MM318 n26 n97 n31 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.205e-05 $Y=0.0001203
MM270 n127 n40 n51 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.995e-05 $Y=0.0001203
MM161 n3 n6 n122 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.415e-05 $Y=4.17e-05
MM111 n73 n8 n110 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.205e-05 $Y=8.85e-05
MM391 n4 Addr1 n62 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001245 $Y=7.35e-05
MM118 n3 n74 n118 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.925e-05 $Y=9.69e-05
MM347 n7 n35 n77 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.945e-05 $Y=1.65e-05
MM358 n4 n66 n22 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.905e-05 $Y=0.0001203
MM120 n3 n106 n76 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.925e-05 $Y=5.01e-05
MM138 n7 n80 n77 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.945e-05 $Y=3.3e-06
MM292 n4 n21 n139 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.945e-05 $Y=0.0001671
MM49 n3 n57 n181 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.245e-05 $Y=4.17e-05
MM258 n4 n57 n181 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.245e-05 $Y=2.67e-05
MM254 n40 n29 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.245e-05 $Y=0.0001203
MM43 n3 n142 n37 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.245e-05 $Y=0.0001821
MM366 n4 n22 n112 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.415e-05 $Y=0.0001203
MM242 n183 n43 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.65e-06 $Y=2.67e-05
MM98 n3 n35 n80 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.455e-05 $Y=3.3e-06
MM132 n153 n131 n72 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.945e-05 $Y=0.0001437
MM184 n3 n147 n161 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001296 $Y=8.85e-05
MM296 n4 n21 n87 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.945e-05 $Y=7.35e-05
MM144 n44 n30 n173 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.185e-05 $Y=5.01e-05
MM114 n20 n80 n151 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.205e-05 $Y=3.3e-06
MM36 n53 n129 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.35e-06 $Y=0.0001437
MM100 n42 n15 n55 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.965e-05 $Y=0.0001437
MM123 n126 n90 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.435e-05 $Y=0.0001821
MM244 n142 n169 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.35e-06 $Y=0.0001671
MM169 n124 n6 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.925e-05 $Y=4.17e-05
MM185 n3 n178 n141 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001347 $Y=9.69e-05
MM11 n174 n93 n160 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.725e-05 $Y=0.0001785
MM279 n4 n146 n98 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.505e-05 $Y=0.0001101
MM222 n103 n93 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.725e-05 $Y=0.0001203
MM332 n126 n90 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.435e-05 $Y=0.0001671
MM350 n112 n59 n66 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.185e-05 $Y=0.0001203
MM218 n43 n96 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.965e-05 $Y=2.67e-05
MM55 n56 n176 n17 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.755e-05 $Y=8.85e-05
MM149 n22 n66 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.905e-05 $Y=0.0001353
MM234 n43 Addr2 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.485e-05 $Y=2.67e-05
MM363 n167 n77 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.905e-05 $Y=1.65e-05
MM103 n73 n87 n113 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.965e-05 $Y=8.85e-05
MM54 n146 n150 n17 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.755e-05 $Y=9.69e-05
MM188 n82 n147 n25 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001419 $Y=8.85e-05
MM45 n40 n29 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.245e-05 $Y=0.0001353
MM414 n107 n101 n177 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001935 $Y=0.0001101
MM400 n166 n178 n65 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001494 $Y=0.0001101
MM134 n118 n99 n164 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.945e-05 $Y=9.69e-05
MM404 n24 n67 n51 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001569 $Y=0.0001101
MM361 n61 n173 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.905e-05 $Y=6.33e-05
MM302 n4 n97 n59 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.455e-05 $Y=0.0001203
MM14 n184 Addr0 n168 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.725e-05 $Y=9.69e-05
MM307 n4 n35 n80 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.455e-05 $Y=1.65e-05
MM95 n3 n87 n8 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.455e-05 $Y=8.85e-05
MM40 n3 n171 n155 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.35e-06 $Y=5.01e-05
MM408 n4 n65 n11 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001665 $Y=0.0001101
MM2 n3 Addr2 n111 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-3.885e-05 $Y=0.0001353
MM171 n154 n149 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.435e-05 $Y=0.0001821
MM381 n52 n158 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.435e-05 $Y=0.0001569
MM108 n42 n131 n86 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.205e-05 $Y=0.0001437
MM416 n105 n177 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000201 $Y=0.0001101
MM107 n152 n46 n126 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.205e-05 $Y=0.0001821
MM182 n3 Addr1 n62 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001245 $Y=8.85e-05
MM51 n17 n37 n144 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.755e-05 $Y=0.0001821
MM239 n4 n33 n157 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.65e-06 $Y=0.0001101
MM22 n33 Addr1 n184 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.485e-05 $Y=9.69e-05
MM16 n148 n93 n180 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.725e-05 $Y=5.01e-05
MM157 n3 n22 n112 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.415e-05 $Y=0.0001353
MM314 n41 n85 n48 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.965e-05 $Y=2.67e-05
MM278 n4 n127 n70 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.505e-05 $Y=0.0001203
MM209 n4 Addr0 n93 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-3.885e-05 $Y=0.0001671
MM84 n3 n21 n15 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.945e-05 $Y=0.0001437
MM286 n38 n70 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.015e-05 $Y=0.0001203
MM135 n125 n8 n92 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.945e-05 $Y=8.85e-05
MM330 n45 n48 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.925e-05 $Y=2.67e-05
MM271 n146 n150 n128 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.995e-05 $Y=0.0001101
MM192 n94 n32 n82 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001494 $Y=8.85e-05
MM194 n94 n62 n172 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001518 $Y=8.85e-05
MM263 n146 n137 n17 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.755e-05 $Y=0.0001101
MM6 n3 n111 n168 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.965e-05 $Y=9.69e-05
MM335 n4 n118 n13 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.435e-05 $Y=0.0001101
MM57 n123 n181 n17 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.755e-05 $Y=4.17e-05
MM326 n4 n26 n159 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.925e-05 $Y=0.0001203
MM275 n78 n145 n89 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.995e-05 $Y=1.65e-05
MM79 n113 n133 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.015e-05 $Y=8.85e-05
MM83 n139 n21 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.945e-05 $Y=0.0001821
MM125 n3 n159 n31 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.435e-05 $Y=0.0001353
MM341 n153 n15 n72 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.945e-05 $Y=0.0001569
MM117 n3 n26 n159 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.925e-05 $Y=0.0001353
MM208 n170 n105 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002061 $Y=9.69e-05
MM373 n158 n115 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.925e-05 $Y=0.0001569
MM264 n56 n120 n17 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.755e-05 $Y=7.35e-05
MM62 n146 n137 n128 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.995e-05 $Y=9.69e-05
MM102 n74 n84 n5 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.965e-05 $Y=9.69e-05
MM3 n174 n96 n3 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.965e-05 $Y=0.0001785
MM213 n4 n111 n16 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.965e-05 $Y=0.0001569
MM71 n3 n56 n133 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.505e-05 $Y=8.85e-05
MM29 n3 n103 n49 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-7.65e-06 $Y=0.0001353
MM405 n50 n147 n172 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001569 $Y=7.35e-05
MM348 n34 n46 n58 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.185e-05 $Y=0.0001671
MM65 n123 n57 n25 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.995e-05 $Y=4.17e-05
MM401 n94 n62 n82 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001494 $Y=7.35e-05
MM86 n3 n21 n84 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.945e-05 $Y=9.69e-05
MM47 n3 n120 n176 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.245e-05 $Y=8.85e-05
MM265 n10 n155 n17 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.755e-05 $Y=6.33e-05
MM93 n3 n97 n59 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.455e-05 $Y=0.0001353
MM324 n90 n152 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.925e-05 $Y=0.0001671
MM24 n180 Addr1 n75 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.485e-05 $Y=5.01e-05
MM410 n4 n11 n54 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001716 $Y=0.0001101
MM247 n4 n157 n137 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.35e-06 $Y=0.0001101
MM146 n143 n35 n77 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.185e-05 $Y=3.3e-06
MM267 n17 n81 n89 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.755e-05 $Y=1.65e-05
MM126 n13 n118 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.435e-05 $Y=9.69e-05
MM160 n44 n61 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.415e-05 $Y=5.01e-05
MM52 n64 n119 n17 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.755e-05 $Y=0.0001437
MM343 n118 n84 n164 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.945e-05 $Y=0.0001101
MM395 n4 n62 n32 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001347 $Y=7.35e-05
MM202 n107 n102 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001716 $Y=8.85e-05
MM121 n3 n48 n45 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.925e-05 $Y=4.17e-05
MM156 n3 n115 n95 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.415e-05 $Y=0.0001437
MM163 n149 n109 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.925e-05 $Y=0.0001821
MM349 n95 n131 n153 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.185e-05 $Y=0.0001569
MM346 n45 n83 n60 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.945e-05 $Y=2.67e-05
MM321 n106 n30 n165 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.205e-05 $Y=6.33e-05
MM284 n162 n23 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.015e-05 $Y=0.0001671
MM245 n4 n129 n53 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.35e-06 $Y=0.0001569
MM9 n9 n96 n3 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.965e-05 $Y=3.81e-05
MM392 n47 n67 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001296 $Y=0.0001101
MM378 n124 n6 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.925e-05 $Y=2.67e-05
MM285 n55 n121 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.015e-05 $Y=0.0001569
MM97 n3 n83 n85 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.455e-05 $Y=4.17e-05
MM375 n88 n39 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.925e-05 $Y=0.0001101
MM417 n170 n105 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002061 $Y=0.0001101
MM110 n74 n99 n13 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.205e-05 $Y=9.69e-05
MM402 n24 n141 n65 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001518 $Y=0.0001101
MM384 n4 n130 n27 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.435e-05 $Y=7.35e-05
MM155 n3 n109 n34 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.415e-05 $Y=0.0001821
MM147 n109 n58 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.905e-05 $Y=0.0001821
MM398 n166 n67 n154 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001443 $Y=0.0001101
MM180 n3 Addr0 n147 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001194 $Y=8.85e-05
MM409 n102 n94 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001665 $Y=7.35e-05
MM272 n56 n176 n27 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.995e-05 $Y=7.35e-05
MM42 n81 n179 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.35e-06 $Y=3.3e-06
MM387 n78 n63 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.435e-05 $Y=1.65e-05
MM38 n137 n157 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.35e-06 $Y=9.69e-05
MM342 n159 n97 n66 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.945e-05 $Y=0.0001203
MM328 n4 n73 n125 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.925e-05 $Y=7.35e-05
MM380 n4 n149 n154 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.435e-05 $Y=0.0001671
MM351 n136 n99 n164 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.185e-05 $Y=0.0001101
MM214 n4 Addr1 n103 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.965e-05 $Y=0.0001203
MM323 n20 n35 n151 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=5.205e-05 $Y=1.65e-05
MM259 n145 n81 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.245e-05 $Y=1.65e-05
MM251 n4 n179 n81 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.35e-06 $Y=1.65e-05
MM129 n28 n45 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.435e-05 $Y=4.17e-05
MM345 n173 n30 n76 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.945e-05 $Y=6.33e-05
MM223 n4 Addr0 n33 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.725e-05 $Y=0.0001101
MM56 n10 n114 n17 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=1.755e-05 $Y=5.01e-05
MM393 n4 n147 n161 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001296 $Y=7.35e-05
MM197 n24 n67 n128 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001593 $Y=9.69e-05
MM88 n3 n21 n30 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.945e-05 $Y=5.01e-05
MM113 n48 n85 n28 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.205e-05 $Y=4.17e-05
MM159 n18 n12 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.415e-05 $Y=8.85e-05
MM81 n41 n36 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=3.015e-05 $Y=4.17e-05
MM411 n107 n102 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001716 $Y=7.35e-05
MM41 n3 n183 n57 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.35e-06 $Y=4.17e-05
MM115 n90 n152 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.925e-05 $Y=0.0001821
MM158 n3 n39 n136 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.415e-05 $Y=9.69e-05
MM277 n121 n64 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.505e-05 $Y=0.0001569
MM151 n12 n92 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.905e-05 $Y=8.85e-05
MM413 n4 n101 n100 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001884 $Y=0.0001101
MM183 n3 n67 n47 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001296 $Y=9.69e-05
MM283 n175 n89 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.505e-05 $Y=1.65e-05
MM200 n102 n94 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001665 $Y=8.85e-05
MM176 n3 n68 n50 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.435e-05 $Y=5.01e-05
MM104 n106 n30 n132 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.965e-05 $Y=5.01e-05
MM288 n4 n133 n113 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.015e-05 $Y=7.35e-05
MM232 n116 Addr2 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.485e-05 $Y=7.35e-05
MM376 n130 n12 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.925e-05 $Y=7.35e-05
MM312 n73 n8 n113 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.965e-05 $Y=7.35e-05
MM23 n117 Addr2 n116 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.485e-05 $Y=8.49e-05
MM1 n3 Addr1 n96 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-3.885e-05 $Y=0.0001437
MM237 n4 n16 n129 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.65e-06 $Y=0.0001569
MM337 n165 n76 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.435e-05 $Y=6.33e-05
MM26 n104 n96 n19 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.485e-05 $Y=3.3e-06
MM69 n3 n127 n70 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.505e-05 $Y=0.0001353
MM74 n175 n89 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.505e-05 $Y=3.3e-06
MM189 n166 n47 n154 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001443 $Y=9.69e-05
MM388 n67 Addr0 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001194 $Y=0.0001101
MM334 n4 n159 n31 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=6.435e-05 $Y=0.0001203
MM274 n123 n181 n25 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.995e-05 $Y=2.67e-05
MM256 n4 n120 n176 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.245e-05 $Y=7.35e-05
MM37 n3 n49 n29 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.35e-06 $Y=0.0001353
MM105 n48 n83 n41 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.965e-05 $Y=4.17e-05
MM253 n119 n53 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.245e-05 $Y=0.0001569
MM224 n4 Addr0 n116 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.725e-05 $Y=7.35e-05
MM371 n4 n167 n143 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.415e-05 $Y=1.65e-05
MM304 n4 n87 n8 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.455e-05 $Y=7.35e-05
MM298 n4 n21 n83 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.945e-05 $Y=2.67e-05
MM216 n4 Addr1 n116 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.965e-05 $Y=7.35e-05
MM206 n54 n101 n177 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001959 $Y=9.69e-05
MM122 n3 n151 n7 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=5.925e-05 $Y=3.3e-06
MM262 n127 n29 n17 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.755e-05 $Y=0.0001203
MM260 n144 n142 n17 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.755e-05 $Y=0.0001671
MM168 n68 n61 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.925e-05 $Y=5.01e-05
MM101 n26 n97 n38 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.965e-05 $Y=0.0001353
MM379 n63 n167 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.925e-05 $Y=1.65e-05
MM294 n4 n21 n97 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.945e-05 $Y=0.0001203
MM293 n15 n21 n4 n4 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=3.945e-05 $Y=0.0001569
MM15 n117 Addr0 n156 n3 C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=-1.725e-05 $Y=8.49e-05
.ENDS
