*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: inv_4x
* View Name: schematic
* Netlist created: 23.Feb.2019 17:45:52
*******************************************************************************

*.SCALE MICRONS
*.GLOBAL vdd gnd

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    inv_4x
* View Name:    schematic
*******************************************************************************

.SUBCKT inv_4x A Z wp=1.6u wn=0.8u lp=0.13u ln=0.13u
*.PININFO Z:O A:I

M1 Z A gnd gnd nch w=3.6 l=0.6 m=2
I5 Z A n1 n1 pch w=7.2 l=0.6 m=2
.ENDS

.END
