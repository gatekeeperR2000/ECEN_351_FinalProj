*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib_bad
* Top Cell Name: or3_1x
* View Name: extracted
* Netlist created: 22.Feb.2025 09:30:50
*******************************************************************************

*.SCALE METER
.GLOBAL vdd
.GLOBAL vss

*******************************************************************************
* Library Name: C5N_std_lib_bad
* Cell Name:    or3_1x
* View Name:    extracted
*******************************************************************************

.SUBCKT or3_1x B Y C A
*.PININFO B:B Y:B C:B A:B

MM10 Y n6 vdd vdd C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.565e-05 $Y=1.53e-05
MM9 vdd A n7 vdd C5NPMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=1.635e-05 $Y=1.35e-05
MM7 n8 C n6 vdd C5NPMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=1.155e-05 $Y=1.35e-05
MM6 n8 C n6 vdd C5NPMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=9.15e-06 $Y=1.35e-05
MM4 vdd A n7 vdd C5NPMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=4.35e-06 $Y=1.35e-05
MM3 Y n6 vss vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.565e-05 $Y=2.1e-06
MM8 n8 B n7 vdd C5NPMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=1.395e-05 $Y=1.35e-05
MM2 vss C n6 vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.15e-06 $Y=2.1e-06
MM1 vss B n6 vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=6.75e-06 $Y=2.1e-06
MM5 n8 B n7 vdd C5NPMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=6.75e-06 $Y=1.35e-05
MM0 vss A n6 vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.35e-06 $Y=2.1e-06
.ENDS
