*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: mux4to1_1x
* View Name: schematic
* Netlist created: 09.Apr.2019 20:36:03
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    mux4to1_1x
* View Name:    schematic
*******************************************************************************

.SUBCKT mux4to1_1x in1 sel1 sel0 in0 in3 out in2 
*.PININFO sel1:I in1:I in0:I sel0:I in2:I out:O in3:I

M29 sel1bb sel1b vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M24 sel1b sel1 vss vss C5NNMOS w=1.8u l=0.6u m=1
M20 mout sel1bb in23 vss C5NNMOS w=1.8u l=0.6u m=1
M2 sel0b sel0 vss vss C5NNMOS w=1.8u l=0.6u m=1
M26 sel1b sel1 vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M26_52 mout sel1bb in01 vdd C5NPMOS w=3.6u l=0.6u m=1
M27 out moutb vss vss C5NNMOS w=1.8u l=0.6u m=1
M22 moutb mout vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M14 in01 sel0b in0 vss C5NNMOS w=1.8u l=0.6u m=1
M0 sel0b sel0 vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M18_46 in23 sel0bb in2 vdd C5NPMOS w=3.6u l=0.6u m=1
M18 moutb mout vss vss C5NNMOS w=1.8u l=0.6u m=1
M17 out moutb vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M28 sel1bb sel1b vss vss C5NNMOS w=1.8u l=0.6u m=1
M23 mout sel1b in23 vdd C5NPMOS w=3.6u l=0.6u m=1
M19 in23 sel0b in2 vss C5NNMOS w=1.8u l=0.6u m=1
M16 in01 sel0bb in1 vss C5NNMOS w=1.8u l=0.6u m=1
M11 in23 sel0b in3 vdd C5NPMOS w=3.6u l=0.6u m=1
M15 in01 sel0b in1 vdd C5NPMOS w=3.6u l=0.6u m=1
M25 mout sel1b in01 vss C5NNMOS w=1.8u l=0.6u m=1
M3 sel0bb sel0b vss vss C5NNMOS w=1.8u l=0.6u m=1
M10_21 in23 sel0bb in3 vss C5NNMOS w=1.8u l=0.6u m=1
M13 in01 sel0bb in0 vdd C5NPMOS w=3.6u l=0.6u m=1
M1 sel0bb sel0b vdd vdd C5NPMOS w=3.6u l=0.6u m=1
.ENDS

