*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: nor2_2x
* View Name: extracted
* Netlist created: 23.Mar.2019 18:06:02
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    nor2_2x
* View Name:    extracted
*******************************************************************************

.SUBCKT nor2_2x Y B
*.PININFO Y:B B:B

MM18 vdd A n5 vdd C5NPMOS w=7.2e-06 l=6e-07 as=5.94e-12 ps=1.77e-05 ad=6.48e-12 pd=1.8e-05 $X=9.15 $Y=11.7
MM14 vss A Y vss C5NNMOS w=1.8e-06 l=6e-07 as=1.485e-12 ps=6.9e-06 ad=1.62e-12 pd=7.2e-06 $X=9.15 $Y=2.1
MM13 Y A vss vss C5NNMOS w=1.8e-06 l=6e-07 as=1.485e-12 ps=6.9e-06 ad=1.62e-12 pd=7.2e-06 $X=6.75 $Y=2.1
MM12 vss B Y vss C5NNMOS w=1.8e-06 l=6e-07 as=1.485e-12 ps=6.9e-06 ad=1.62e-12 pd=7.2e-06 $X=4.35 $Y=2.1
MM19 n5 B Y vdd C5NPMOS w=7.2e-06 l=6e-07 as=5.94e-12 ps=1.77e-05 ad=6.48e-12 pd=1.8e-05 $X=11.55 $Y=11.7
MM17 n5 A vdd vdd C5NPMOS w=7.2e-06 l=6e-07 as=5.94e-12 ps=1.77e-05 ad=6.48e-12 pd=1.8e-05 $X=6.75 $Y=11.7
MM16 Y B n5 vdd C5NPMOS w=7.2e-06 l=6e-07 as=5.94e-12 ps=1.77e-05 ad=6.48e-12 pd=1.8e-05 $X=4.35 $Y=11.7
MM15 Y B vss vss C5NNMOS w=1.8e-06 l=6e-07 as=1.485e-12 ps=6.9e-06 ad=1.62e-12 pd=7.2e-06 $X=11.55 $Y=2.1
.ENDS
