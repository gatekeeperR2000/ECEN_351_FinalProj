*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib_bad
* Top Cell Name: nand2_1x
* View Name: schematic
* Netlist created: 22.Feb.2025 10:42:40
*******************************************************************************

*.SCALE METER
.GLOBAL vdd
.GLOBAL vss

*******************************************************************************
* Library Name: C5N_std_lib_bad
* Cell Name:    nand2_1x
* View Name:    schematic
*******************************************************************************

.SUBCKT nand2_1x B Y A 
*.PININFO Y:O B:I A:I

M3 Y B vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M1 Y A n0 vss C5NNMOS w=3.6u l=0.6u m=1
M2 n0 B vss vss C5NNMOS w=3.6u l=0.6u m=1
M0 Y A vdd vdd C5NPMOS w=3.6u l=0.6u m=1
.ENDS

