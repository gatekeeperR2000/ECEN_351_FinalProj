*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: nand2_4x
* View Name: schematic
* Netlist created: 28.Mar.2019 17:11:57
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    nand2_4x
* View Name:    schematic
*******************************************************************************

.SUBCKT nand2_4x B Y A 
*.PININFO B:I Y:O A:I

M3 Y B vdd vdd C5NPMOS w=3.6u l=0.6u m=4
M1 Y A n0 vss C5NNMOS w=3.6u l=0.6u m=4
M2 n0 B vss vss C5NNMOS w=3.6u l=0.6u m=4
M0 Y A vdd vdd C5NPMOS w=3.6u l=0.6u m=4
.ENDS

