*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: nand3_1x
* View Name: extracted
* Netlist created: 22.Mar.2019 21:21:24
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    nand3_1x
* View Name:    extracted
*******************************************************************************

.SUBCKT nand3_1x Y B C A
*.PININFO Y:B B:B C:B A:B

MM84 Y B vdd vdd C5NPMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=6.75 $Y=15.3
MM81 n6 B n7 vss C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=6.75 $Y=2.1
MM85 vdd A Y vdd C5NPMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=9.15 $Y=15.3
MM83 vdd C Y vdd C5NPMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=4.35 $Y=15.3
MM82 n7 A Y vss C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=9.15 $Y=2.1
MM80 vss C n6 vss C5NNMOS w=5.4e-06 l=6e-07 as=4.455e-12 ps=1.41e-05 ad=4.86e-12 pd=1.44e-05 $X=4.35 $Y=2.1
.ENDS
