* C:\Users\Randall_Jack\Desktop\glade5_win64\ECEN351\C5N_LTspice\buffer_top.asc
XX1 IN OUT POS NEG buffer
V1 NEG 0 0
V2 POS 0 5
V3 IN 0 PULSE(0 5 0 .1n .1n 0.4n 1n)

* block symbol definitions
.subckt buffer IN OUT POS NEG
XX1 IN N001 POS NEG inverter
XX2 N001 OUT POS NEG inverter
.ends buffer

.subckt inverter Vin Vout Vpos Vneg
M1 Vout Vin Vpos Vpos C5NPMOS l=0.6u w=1.8u
M2 Vout Vin Vneg Vneg C5NNMOS l=0.6u w=3.6u
.ends inverter

.model NMOS NMOS
.model PMOS PMOS
.lib C:\Users\Randall_Jack\Documents\LTspiceXVII\lib\cmp\standard.mos
.tran 5n
.include "C5N_models_Glade.txt"
.backanno
.end
