*******************************************************************************
* CDL netlist
*
* Library : buffer_ex
* Top Cell Name: inverter
* View Name: schematic
* Netlist created: 23.Feb.2019 15:57:18
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd gnd

*******************************************************************************
* Library Name: buffer_ex
* Cell Name:    inverter
* View Name:    schematic
*******************************************************************************

.SUBCKT inverter Vin vpos vneg Vout
*.PININFO Vin:I vpos:B Vout:O vneg:B

M1 Vout Vin vneg vneg nch w=1.8u l=0.6u m=1
M0 Vout Vin vpos vpos pch w=1.8u l=0.6u m=1
.ENDS

.END
