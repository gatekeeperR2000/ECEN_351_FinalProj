*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: mux4to1_1x
* View Name: layout
* Netlist created: 09.Apr.2019 20:35:20
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    mux4to1_1x
* View Name:    layout
*******************************************************************************

.SUBCKT mux4to1_1x

.ENDS
