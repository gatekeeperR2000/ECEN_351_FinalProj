*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: mux2to1_1x
* View Name: extracted
* Netlist created: 09.Apr.2019 21:37:41
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    mux2to1_1x
* View Name:    extracted
*******************************************************************************

.SUBCKT mux2to1_1x in1 sel in0 out
*.PININFO in1:B sel:B in0:B out:B

MM20 in1 selb n8 vdd C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=14.55 $Y=15.3
MM13 vss selb selbb vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.45 $Y=2.1
MM15 n8 selb in0 vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=16.95 $Y=2.1
MM14 in1 selbb n8 vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=14.55 $Y=2.1
MM21 n8 selbb in0 vdd C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=16.95 $Y=15.3
MM17 vss n9 out vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=27.15 $Y=2.1
MM19 vdd selb selbb vdd C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.45 $Y=15.3
MM22 vdd n8 n9 vdd C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=22.05 $Y=15.3
MM18 vdd sel selb vdd C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=4.35 $Y=15.3
MM16 vss n8 n9 vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=22.05 $Y=2.1
MM12 vss sel selb vss C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=4.35 $Y=2.1
MM23 vdd n9 out vdd C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=27.15 $Y=15.3
.ENDS
