*******************************************************************************
* CDL netlist
*
* Library : Amplifier
* Top Cell Name: diffamp
* View Name: extracted
* Netlist created: 21.Mar.2019 10:08:32
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: Amplifier
* Cell Name:    diffamp
* View Name:    extracted
*******************************************************************************

.SUBCKT diffamp gnd vinp ibias vinn vout
*.PININFO gnd:B vinp:B ibias:B vinn:B vout:B

MM9 gnd vinn vout gnd C5NNMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=45.9 $Y=15.3
MM6 vout vinn gnd gnd C5NNMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=34.2 $Y=15.3
MM4 n6 vinp gnd gnd C5NNMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=26.4 $Y=15.3
MM7 gnd vinp n6 gnd C5NNMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=38.1 $Y=15.3
MM5 gnd vinn vout gnd C5NNMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=30.3 $Y=15.3
MM2 gnd ibias n7 gnd C5NNMOS w=9.9e-06 l=1.2e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=14.7 $Y=15.3
MM13 vdd n6 vout vdd C5NPMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=30.3 $Y=31.35
MM8 n6 vinp gnd gnd C5NNMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=42 $Y=15.3
MM3 gnd vinp n6 gnd C5NNMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=22.5 $Y=15.3
MM15 vdd n6 n6 vdd C5NPMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=38.1 $Y=31.35
MM14 vout n6 vdd vdd C5NPMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=34.2 $Y=31.35
MM17 vdd n6 vout vdd C5NPMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=45.9 $Y=31.35
MM18 vout n6 vdd vdd C5NPMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=49.8 $Y=31.35
MM16 n6 n6 vdd vdd C5NPMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=42 $Y=31.35
MM12 n6 n6 vdd vdd C5NPMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=26.4 $Y=31.35
MM10 vout vinn gnd gnd C5NNMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=49.8 $Y=15.3
MM11 vdd n6 n6 vdd C5NPMOS w=9.9e-06 l=2.1e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=22.5 $Y=31.35
MM0 ibias ibias gnd gnd C5NNMOS w=9.9e-06 l=1.2e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=8.7 $Y=15.3
MM1 gnd ibias gnd gnd C5NNMOS w=9.9e-06 l=1.2e-06 as=1.6335e-11 ps=2.31e-05 ad=1.782e-11 pd=2.34e-05 $X=11.7 $Y=15.3
.ENDS
