*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: mux2to1_1x
* View Name: schematic
* Netlist created: 09.Apr.2019 21:37:40
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    mux2to1_1x
* View Name:    schematic
*******************************************************************************

.SUBCKT mux2to1_1x sel in1 in0 out 
*.PININFO sel:I in1:I in0:I out:O

M9 n6 n2 vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M10_21 n2 selbb in1 vss C5NNMOS w=1.8u l=0.6u m=1
M2 selb sel vss vss C5NNMOS w=1.8u l=0.6u m=1
M8 n6 n2 vss vss C5NNMOS w=1.8u l=0.6u m=1
M3 selbb selb vss vss C5NNMOS w=1.8u l=0.6u m=1
M18 n2 selbb in0 vdd C5NPMOS w=3.6u l=0.6u m=1
M19 n2 selb in0 vss C5NNMOS w=1.8u l=0.6u m=1
M12 out n6 vss vss C5NNMOS w=1.8u l=0.6u m=1
M10 out n6 vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M11 n2 selb in1 vdd C5NPMOS w=3.6u l=0.6u m=1
M0 selb sel vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M1 selbb selb vdd vdd C5NPMOS w=3.6u l=0.6u m=1
.ENDS

