*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: inv_8x
* View Name: schematic
* Netlist created: 22.Mar.2019 20:49:56
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    inv_8x
* View Name:    schematic
*******************************************************************************

.SUBCKT inv_8x Z A 
*.PININFO Z:O A:I

M4 Z A vss vss C5NNMOS w=1.8u l=0.6u m=8
M5 Z A vdd vdd C5NPMOS w=3.6u l=0.6u m=8
.ENDS

