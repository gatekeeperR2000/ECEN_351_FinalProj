*******************************************************************************
* CDL netlist
*
* Library : buffer_ex
* Top Cell Name: inverter
* View Name: schematic
* Netlist created: 23.Feb.2019 20:53:21
*******************************************************************************

*.SCALE MICRONS
*.GLOBAL vpos vneg

*******************************************************************************
* Library Name: buffer_ex
* Cell Name:    inverter
* View Name:    schematic
*******************************************************************************

.SUBCKT inverter Vin Vout
*.PININFO Vout:O Vin:I

M0 Vout Vin vpos vpos pch
M1 vneg vneg Vout Vin nch
.ENDS

