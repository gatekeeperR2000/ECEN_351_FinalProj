*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: nor3_1x
* View Name: schematic
* Netlist created: 31.Aug.2023 15:08:28
*******************************************************************************

*.SCALE METER
.GLOBAL vdd
.GLOBAL vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    nor3_1x
* View Name:    schematic
*******************************************************************************

.SUBCKT nor3_1x B Y A 
*.PININFO B:I Y:O C:I A:I

M4 Y C vss vss C5NNMOS w=1.8u l=0.6u m=1
M2 Y B vss vss C5NNMOS w=1.8u l=0.6u m=1
M5 Y C n2 vdd C5NPMOS w=10.8u l=0.6u m=1
M3 n2 B n3 vdd C5NPMOS w=10.8u l=0.6u m=1
M1 Y A vss vss C5NNMOS w=1.8u l=0.6u m=1
M0 n3 A vdd vdd C5NPMOS w=10.8u l=0.6u m=1
.ENDS

