*******************************************************************************
* CDL netlist
*
* Library : buffer_ex
* Top Cell Name: inverter
* View Name: schematic
* Netlist created: 23.Feb.2019 22:44:16
*******************************************************************************

*.SCALE METER
*.GLOBAL vpos vneg

*******************************************************************************
* Library Name: buffer_ex
* Cell Name:    inverter
* View Name:    schematic
*******************************************************************************

.SUBCKT inverter Vin Vout
*.PININFO Vout:O Vin:I

M1 Vout Vin vneg vneg C5NNMOS w=1.8u l=0.6u m=1
M0 Vout Vin vpos vpos C5NPMOS w=1.8u l=0.6u m=1
.ENDS

