*******************************************************************************
* CDL netlist
*
* Library : buffer_ex
* Top Cell Name: inverter
* View Name: schematic
* Netlist created: 23.Feb.2019 21:20:57
*******************************************************************************

*.SCALE METER
*.GLOBAL vpos vneg

*******************************************************************************
* Library Name: buffer_ex
* Cell Name:    inverter
* View Name:    schematic
*******************************************************************************

.SUBCKT inverter Vin Vout
*.PININFO Vin:I Vout:O

M1 Vin Vout vneg vneg nch
M0 vpos vpos Vin Vout pch
.ENDS

.END
