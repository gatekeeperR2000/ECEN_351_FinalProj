*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: D_Flip_Flop
* View Name: schematic
* Netlist created: 04.Mar.2025 07:57:06
*******************************************************************************

*.SCALE METER
.GLOBAL vdd
.GLOBAL vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    D_Flip_Flop
* View Name:    schematic
*******************************************************************************

.SUBCKT D_Flip_Flop D_in clk Q_out Qn_out 
*.PININFO D_in:I Q_out:O clk:I Qn_out:O

M20 n15 n11 vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M2 clkb clk vss vss C5NNMOS w=1.8u l=0.6u m=1
M22 n6 clkbb n11 vdd C5NPMOS w=3.6u l=0.6u m=1
M14 n3 n12 vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M0 clkb clk vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M12 n3 clkb n9 vdd C5NPMOS w=3.6u l=0.6u m=1
M4 Q_out Qn_out vss vss C5NNMOS w=1.8u l=0.6u m=1
M6 Qn_out n15 vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M18 n11 clkb n12 vdd C5NPMOS w=3.6u l=0.6u m=1
M17 n6 clkb n11 vss C5NNMOS w=1.8u l=0.6u m=1
M23 n6 n15 vss vss C5NNMOS w=1.8u l=0.6u m=1
M19 n11 clkbb n12 vss C5NNMOS w=1.8u l=0.6u m=1
M9 n12 n9 vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M11 n9 clkbb D_in vdd C5NPMOS w=3.6u l=0.6u m=1
M16 n6 n15 vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M15 n3 n12 vss vss C5NNMOS w=1.8u l=0.6u m=1
M5 Q_out Qn_out vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M21 n15 n11 vss vss C5NNMOS w=1.8u l=0.6u m=1
M3 clkbb clkb vss vss C5NNMOS w=1.8u l=0.6u m=1
M7 Qn_out n15 vss vss C5NNMOS w=1.8u l=0.6u m=1
M8 n12 n9 vss vss C5NNMOS w=1.8u l=0.6u m=1
M13 n3 clkbb n9 vss C5NNMOS w=1.8u l=0.6u m=1
M1 clkbb clkb vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M10 n9 clkb D_in vss C5NNMOS w=1.8u l=0.6u m=1
.ENDS

.END
