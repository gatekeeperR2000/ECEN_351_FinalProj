*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: and2_4x
* View Name: schematic
* Netlist created: 22.Mar.2019 20:11:26
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    and2_4x
* View Name:    schematic
*******************************************************************************

.SUBCKT and2_4x B Y A 
*.PININFO B:I Y:O A:I

M4 Y n0 vss vss C5NNMOS w=1.8u l=0.6u m=4
M2 n2 B vss vss C5NNMOS w=3.6u l=0.6u m=1
M5 Y n0 vdd vdd C5NPMOS w=3.6u l=0.6u m=4
M3 n0 B vdd vdd C5NPMOS w=3.6u l=0.6u m=1
M1 n0 A n2 vss C5NNMOS w=3.6u l=0.6u m=1
M0 n0 A vdd vdd C5NPMOS w=3.6u l=0.6u m=1
.ENDS

