*******************************************************************************
* CDL netlist
*
* Library : final_version
* Top Cell Name: final_layout
* View Name: extracted
* Netlist created: 03.Apr.2023 13:21:43
*******************************************************************************

*.SCALE METER
.GLOBAL vdd
.GLOBAL vss

*******************************************************************************
* Library Name: final_version
* Cell Name:    final_layout
* View Name:    extracted
*******************************************************************************

.SUBCKT final_layout

MM1200 n83 n5 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-4.83e-05 $Y=-4.17e-05
MM1035 n112 n173 n156 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.46e-05 $Y=-0.00011445
MM1304 n164 n105 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001092 $Y=-0.00013185
MM1318 n108 n179 n71 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001167 $Y=-7.08e-05
MM1369 n6 n163 n111 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001488 $Y=-0.00016245
MM1307 n98 n16 n209 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001143 $Y=2.055e-05
MM1058 n179 n197 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001041 $Y=-8.4e-05
MM1045 n3 n40 n171 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.97e-05 $Y=-0.00017565
MM953 n219 n97 n79 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-8.175e-05 $Y=-6.54e-05
MM950 n89 n165 n166 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-8.415e-05 $Y=-5.49e-05
MM949 n3 n86 n178 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-9.135e-05 $Y=-6.18e-05
MM1096 n3 n134 n194 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000129 $Y=-2.235e-05
MM960 n205 n97 n1 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-6.03e-05 $Y=-5.49e-05
MM1170 n158 n138 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002595 $Y=-5.49e-05
MM1359 n31 n99 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001437 $Y=-0.00010125
MM1196 n130 n97 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-6.03e-05 $Y=-4.17e-05
MM1099 n126 n18 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000129 $Y=-0.00011445
MM1383 n6 n84 n112 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000159 $Y=-0.00010125
MM1267 n36 n203 n24 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.46e-05 $Y=2.055e-05
MM1362 n6 n106 n91 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001488 $Y=5.1e-05
MM955 n3 n41 n79 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-7.935e-05 $Y=-6.54e-05
MM1159 n182 n2 n24 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00023505 $Y=-3.93e-05
MM990 n159 n22 n66 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=2.175e-05 $Y=3.78e-05
MM967 n52 n165 n141 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-4.11e-05 $Y=-6.54e-05
MM952 n217 n97 n166 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-8.175e-05 $Y=-5.49e-05
MM1116 n151 n105 n78 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001365 $Y=-0.00014505
MM1103 n72 n16 n29 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001341 $Y=7.35e-06
MM944 n11 n165 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=-0.00010335 $Y=-5.49e-05
MM1410 n109 n81 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00029415 $Y=-3.735e-05
MM1343 n99 n30 n18 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001341 $Y=-0.00010125
MM997 n225 n178 n162 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=2.175e-05 $Y=-0.00017565
MM1370 n170 n106 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001539 $Y=5.1e-05
MM1174 n3 n81 n109 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00029415 $Y=-5.055e-05
MM1306 n174 n26 n44 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001143 $Y=5.1e-05
MM1034 n20 n120 n149 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.46e-05 $Y=-8.4e-05
MM1405 n58 n118 n125 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00025245 $Y=-2.61e-05
MM1056 n45 n198 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001041 $Y=-2.235e-05
MM1312 n107 n164 n132 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001143 $Y=-0.00013185
MM1081 n147 n85 n161 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001167 $Y=-5.355e-05
MM1121 n95 n28 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001437 $Y=-5.355e-05
MM1141 n19 n163 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001539 $Y=-0.00017565
MM1268 n68 n93 n27 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.46e-05 $Y=-9.15e-06
MM1319 n208 n30 n126 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001167 $Y=-0.00010125
MM1005 n3 n162 n139 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.895e-05 $Y=-0.00017565
MM1154 n3 n145 n115 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002226 $Y=-5.49e-05
MM1049 n92 n154 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.48e-05 $Y=-5.355e-05
MM1079 n98 n16 n13 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001167 $Y=7.35e-06
MM1230 n103 n62 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.175e-05 $Y=-7.08e-05
MM1024 n12 n93 n27 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.22e-05 $Y=-2.235e-05
MM1142 n3 n170 n188 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000159 $Y=3.78e-05
MM988 n223 n144 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=1.935e-05 $Y=-0.00014505
MM1199 n6 n41 n129 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-5.79e-05 $Y=-7.68e-05
MM1063 n3 n4 n16 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001092 $Y=7.35e-06
MM978 n3 n54 n221 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-1.47e-05 $Y=-5.49e-05
MM1315 n98 n4 n13 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001167 $Y=2.055e-05
MM1131 n3 n31 n37 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001488 $Y=-0.00011445
MM1015 n3 n80 n203 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.71e-05 $Y=7.35e-06
MM980 n41 n54 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=-3e-06 $Y=-5.49e-05
MM966 n5 n165 n153 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-4.11e-05 $Y=-5.49e-05
MM1387 n6 n119 n2 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00021255 $Y=-2.61e-05
MM959 n129 n11 n122 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-6.27e-05 $Y=-6.54e-05
MM1105 n90 n85 n28 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001341 $Y=-5.355e-05
MM1272 n175 n82 n124 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.46e-05 $Y=-0.00013185
MM1339 n72 n4 n29 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001341 $Y=2.055e-05
MM1195 n6 n11 n129 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-6.27e-05 $Y=-7.68e-05
MM1303 n6 n30 n38 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001092 $Y=-0.00010125
MM1155 n118 n2 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00022275 $Y=-3.93e-05
MM1349 n74 n85 n28 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001365 $Y=-4.035e-05
MM969 n210 n113 n141 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-3.87e-05 $Y=-6.54e-05
MM1201 n6 n52 n123 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-4.83e-05 $Y=-7.68e-05
MM1249 n10 n139 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.2e-05 $Y=-0.00016245
MM1120 n3 n76 n167 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001437 $Y=-2.235e-05
MM1158 n192 n145 n124 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002349 $Y=-5.49e-05
MM1090 n3 n108 n146 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001239 $Y=-8.4e-05
MM1108 n150 n164 n78 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001341 $Y=-0.00014505
MM1083 n208 n38 n126 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001167 $Y=-0.00011445
MM1382 n20 n53 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000159 $Y=-7.08e-05
MM1403 n68 n2 n125 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00025005 $Y=-2.61e-05
MM1156 n3 n196 n117 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002277 $Y=-5.49e-05
MM965 n3 n52 n123 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-4.83e-05 $Y=-6.18e-05
MM1391 n6 n2 n118 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00022275 $Y=-2.61e-05
MM1214 n33 n54 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.47e-05 $Y=-4.17e-05
MM1337 n195 n0 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000129 $Y=-0.00016245
MM1309 n147 n85 n140 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001143 $Y=-4.035e-05
MM1091 n3 n208 n18 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001239 $Y=-0.00011445
MM1047 n70 n9 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.48e-05 $Y=7.35e-06
MM1393 n6 n7 n177 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00022785 $Y=-2.61e-05
MM1346 n91 n26 n8 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001365 $Y=5.1e-05
MM1071 n98 n4 n209 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001143 $Y=7.35e-06
MM1353 n111 n191 n64 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001365 $Y=-0.00016245
MM1133 n111 n163 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001488 $Y=-0.00017565
MM963 n3 n41 n226 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-5.79e-05 $Y=-6.54e-05
MM1014 n3 n15 n180 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.71e-05 $Y=3.78e-05
MM1367 n37 n31 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001488 $Y=-0.00010125
MM1372 n47 n167 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001539 $Y=-9.15e-06
MM1019 n3 n173 n46 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.71e-05 $Y=-0.00011445
MM1380 n6 n47 n68 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000159 $Y=-9.15e-06
MM1114 n193 n179 n148 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001365 $Y=-8.4e-05
MM1298 n6 n121 n26 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001092 $Y=5.1e-05
MM1017 n184 n96 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.71e-05 $Y=-5.355e-05
MM1245 n96 n183 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.2e-05 $Y=-4.035e-05
MM999 n135 n137 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.895e-05 $Y=7.35e-06
MM1357 n6 n28 n95 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001437 $Y=-4.035e-05
MM986 n3 n144 n201 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=1.935e-05 $Y=-8.4e-05
MM1285 n92 n154 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.48e-05 $Y=-4.035e-05
MM1032 n68 n51 n27 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.46e-05 $Y=-2.235e-05
MM1238 n6 n103 n55 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.895e-05 $Y=-7.08e-05
MM1259 n12 n80 n36 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.22e-05 $Y=2.055e-05
MM1397 n188 n2 n182 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00023745 $Y=-2.61e-05
MM1216 n41 n54 n6 n6 C5NPMOS w=7.2e-06 l=6e-07 as=1.296e-11 ps=1.8e-05 ad=1.188e-11 pd=1.77e-05 $X=-3e-06 $Y=-4.53e-05
MM968 n127 n113 n153 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-3.87e-05 $Y=-5.49e-05
MM1274 n87 n67 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.97e-05 $Y=5.1e-05
MM1246 n6 n55 n120 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.2e-05 $Y=-7.08e-05
MM1179 n60 n25 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00031695 $Y=-5.055e-05
MM1341 n90 n77 n28 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001341 $Y=-4.035e-05
MM1188 n89 n97 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-8.175e-05 $Y=-4.17e-05
MM1404 n20 n115 n102 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002523 $Y=-6.99e-05
MM1352 n151 n164 n78 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001365 $Y=-0.00013185
MM1109 n0 n191 n64 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001341 $Y=-0.00017565
MM1250 n6 n15 n180 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.71e-05 $Y=5.1e-05
MM1051 n73 n104 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.48e-05 $Y=-0.00011445
MM1223 n39 n144 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.935e-05 $Y=-0.00010125
MM1172 n131 n158 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002646 $Y=-5.49e-05
MM1065 n3 n77 n85 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001092 $Y=-5.355e-05
MM1210 n33 n11 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.95e-05 $Y=-4.17e-05
MM1261 n12 n96 n50 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.22e-05 $Y=-4.035e-05
MM1046 n187 n87 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.48e-05 $Y=3.78e-05
MM1016 n3 n51 n93 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.71e-05 $Y=-2.235e-05
MM1018 n3 n120 n181 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.71e-05 $Y=-8.4e-05
MM951 n219 n165 n86 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-8.415e-05 $Y=-6.54e-05
MM1167 n125 n118 n68 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00025005 $Y=-3.93e-05
MM1042 n186 n149 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.97e-05 $Y=-8.4e-05
MM985 n3 n144 n215 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=1.935e-05 $Y=-5.355e-05
MM1409 n23 n189 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00026475 $Y=-2.61e-05
MM1007 n80 n135 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.2e-05 $Y=7.35e-06
MM971 n210 n41 n3 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-3.63e-05 $Y=-6.54e-05
MM1244 n51 n35 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.2e-05 $Y=-9.15e-06
MM1064 n3 n45 n213 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001092 $Y=-2.235e-05
MM1069 n191 n136 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001092 $Y=-0.00017565
MM1347 n63 n16 n72 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001365 $Y=2.055e-05
MM1251 n6 n80 n203 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.71e-05 $Y=2.055e-05
MM1211 n6 n11 n14 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.95e-05 $Y=-7.68e-05
MM1358 n200 n148 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001437 $Y=-7.08e-05
MM1118 n3 n8 n106 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001437 $Y=3.78e-05
MM1310 n108 n204 n49 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001143 $Y=-7.08e-05
MM1030 n188 n15 n67 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.46e-05 $Y=3.78e-05
MM1263 n156 n173 n12 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.22e-05 $Y=-0.00010125
MM1080 n59 n213 n194 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001167 $Y=-2.235e-05
MM1198 n130 n54 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-5.79e-05 $Y=-4.17e-05
MM1057 n77 n199 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001041 $Y=-5.355e-05
MM1281 n171 n40 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.97e-05 $Y=-0.00016245
MM1378 n188 n170 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000159 $Y=5.1e-05
MM1048 n61 n211 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.48e-05 $Y=-2.235e-05
MM1025 n50 n184 n12 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.22e-05 $Y=-5.355e-05
MM1012 n114 n160 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.2e-05 $Y=-0.00014505
MM1224 n185 n144 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.935e-05 $Y=-0.00013185
MM1220 n6 n144 n57 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.935e-05 $Y=-9.15e-06
MM1088 n3 n59 n134 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001239 $Y=-2.235e-05
MM1060 n105 n157 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001041 $Y=-0.00014505
MM1068 n3 n105 n164 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001092 $Y=-0.00014505
MM1143 n24 n142 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000159 $Y=7.35e-06
MM1183 n6 n97 n113 n6 C5NPMOS w=7.2e-06 l=6e-07 as=1.296e-11 ps=1.8e-05 ad=1.188e-11 pd=1.77e-05 $X=-0.00010095 $Y=-7.68e-05
MM946 n11 n165 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=-0.00010095 $Y=-5.49e-05
MM1398 n138 n196 n192 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002424 $Y=-6.99e-05
MM1284 n61 n211 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.48e-05 $Y=-9.15e-06
MM1115 n37 n30 n99 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001365 $Y=-0.00011445
MM1070 n174 n121 n44 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001143 $Y=3.78e-05
MM989 n225 n144 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=1.935e-05 $Y=-0.00017565
MM1368 n6 n169 n151 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001488 $Y=-0.00013185
MM1371 n142 n65 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001539 $Y=2.055e-05
MM1231 n39 n123 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.175e-05 $Y=-0.00010125
MM1008 n51 n35 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.2e-05 $Y=-2.235e-05
MM1122 n200 n148 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001437 $Y=-8.4e-05
MM1269 n58 n184 n50 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.46e-05 $Y=-4.035e-05
MM1001 n183 n94 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.895e-05 $Y=-5.355e-05
MM973 n62 n14 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-2.67e-05 $Y=-6.18e-05
MM1356 n167 n76 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001437 $Y=-9.15e-06
MM1110 n91 n121 n8 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001365 $Y=3.78e-05
MM1150 n3 n119 n145 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002124 $Y=-5.49e-05
MM1127 n3 n65 n63 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001488 $Y=7.35e-06
MM1003 n133 n39 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.895e-05 $Y=-0.00011445
MM1260 n12 n51 n27 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.22e-05 $Y=-9.15e-06
MM1348 n76 n213 n43 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001365 $Y=-9.15e-06
MM1336 n56 n150 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000129 $Y=-0.00013185
MM1209 n6 n14 n62 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-2.67e-05 $Y=-7.68e-05
MM1077 n69 n136 n143 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001143 $Y=-0.00017565
MM1266 n188 n180 n67 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.46e-05 $Y=5.1e-05
MM1322 n32 n174 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001239 $Y=5.1e-05
MM982 n66 n144 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=1.935e-05 $Y=3.78e-05
MM1194 n130 n11 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-6.27e-05 $Y=-4.17e-05
MM1333 n6 n90 n161 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000129 $Y=-4.035e-05
MM983 n101 n144 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=1.935e-05 $Y=7.35e-06
MM1396 n116 n145 n192 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002373 $Y=-6.99e-05
MM962 n3 n54 n1 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-5.79e-05 $Y=-5.49e-05
MM1305 n6 n136 n191 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001092 $Y=-0.00016245
MM1365 n74 n95 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001488 $Y=-4.035e-05
MM1097 n161 n90 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000129 $Y=-5.355e-05
MM1125 n163 n64 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001437 $Y=-0.00017565
MM1162 n138 n117 n192 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002424 $Y=-5.49e-05
MM1308 n59 n213 n88 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001143 $Y=-9.15e-06
MM1233 n162 n178 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.175e-05 $Y=-0.00016245
MM1377 n6 n163 n19 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001539 $Y=-0.00016245
MM1002 n55 n103 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.895e-05 $Y=-8.4e-05
MM1129 n3 n95 n74 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001488 $Y=-5.355e-05
MM1229 n6 n206 n94 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.175e-05 $Y=-4.035e-05
MM1160 n116 n115 n192 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002373 $Y=-5.49e-05
MM1052 n172 n216 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.48e-05 $Y=-0.00014505
MM964 n83 n5 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-4.83e-05 $Y=-5.49e-05
MM961 n122 n97 n226 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-6.03e-05 $Y=-6.54e-05
MM1013 n10 n139 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.2e-05 $Y=-0.00017565
MM1004 n160 n185 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.895e-05 $Y=-0.00014505
MM1027 n156 n46 n12 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.22e-05 $Y=-0.00011445
MM1126 n3 n106 n91 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001488 $Y=3.78e-05
MM1033 n58 n96 n50 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.46e-05 $Y=-5.355e-05
MM1286 n6 n186 n34 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.48e-05 $Y=-7.08e-05
MM1136 n47 n167 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001539 $Y=-2.235e-05
MM1075 n208 n30 n176 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001143 $Y=-0.00011445
MM1100 n56 n150 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000129 $Y=-0.00014505
MM1237 n183 n94 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.895e-05 $Y=-4.035e-05
MM1289 n6 n171 n143 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.48e-05 $Y=-0.00016245
MM1020 n82 n114 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.71e-05 $Y=-0.00014505
MM1006 n3 n42 n15 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.2e-05 $Y=3.78e-05
MM1292 n45 n198 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001041 $Y=-9.15e-06
MM995 n128 n123 n39 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=2.175e-05 $Y=-0.00011445
MM1189 n86 n97 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-8.175e-05 $Y=-7.68e-05
MM1092 n150 n107 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001239 $Y=-0.00014505
MM1363 n6 n65 n63 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001488 $Y=2.055e-05
MM1218 n159 n144 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.935e-05 $Y=5.1e-05
MM1415 n6 n25 n60 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00031695 $Y=-3.735e-05
MM1340 n134 n45 n76 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001341 $Y=-9.15e-06
MM1219 n6 n144 n137 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.935e-05 $Y=2.055e-05
MM1067 n38 n30 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001092 $Y=-0.00011445
MM1270 n149 n181 n20 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.46e-05 $Y=-7.08e-05
MM1178 n25 n100 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00031185 $Y=-5.055e-05
MM1192 n17 n130 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-6.99e-05 $Y=-4.17e-05
MM1175 n3 n109 n21 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00029925 $Y=-5.055e-05
MM1271 n112 n46 n156 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.46e-05 $Y=-0.00010125
MM1152 n3 n75 n196 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002175 $Y=-5.49e-05
MM1278 n6 n149 n186 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.97e-05 $Y=-7.08e-05
MM1193 n6 n129 n207 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-6.99e-05 $Y=-7.68e-05
MM1078 n174 n26 n152 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001167 $Y=3.78e-05
MM1332 n6 n134 n194 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000129 $Y=-9.15e-06
MM1399 n48 n7 n182 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00024255 $Y=-2.61e-05
MM1392 n117 n196 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002277 $Y=-6.99e-05
MM992 n218 n17 n57 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=2.175e-05 $Y=-2.235e-05
MM1389 n6 n75 n7 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00021765 $Y=-2.61e-05
MM1412 n100 n109 n131 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00030435 $Y=-3.735e-05
MM1360 n169 n78 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001437 $Y=-0.00013185
MM1381 n58 n212 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000159 $Y=-4.035e-05
MM1106 n148 n204 n146 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001341 $Y=-8.4e-05
MM1191 n6 n41 n86 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.935e-05 $Y=-7.68e-05
MM1243 n80 n135 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.2e-05 $Y=2.055e-05
MM1168 n20 n145 n102 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002523 $Y=-5.49e-05
MM996 n223 n207 n185 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=2.175e-05 $Y=-0.00014505
MM1330 n152 n32 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000129 $Y=5.1e-05
MM1320 n107 n105 n56 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001167 $Y=-0.00013185
MM1208 n22 n33 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-2.67e-05 $Y=-4.17e-05
MM1197 n6 n97 n129 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-6.03e-05 $Y=-7.68e-05
MM976 n202 n113 n221 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-1.71e-05 $Y=-5.49e-05
MM947 n3 n97 n113 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=-0.00010095 $Y=-6.36e-05
MM1145 n3 n212 n58 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000159 $Y=-5.355e-05
MM1132 n151 n169 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001488 $Y=-0.00014505
MM1277 n154 n50 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.97e-05 $Y=-4.035e-05
MM1240 n160 n185 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.895e-05 $Y=-0.00013185
MM991 n101 n83 n137 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=2.175e-05 $Y=7.35e-06
MM1296 n105 n157 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001041 $Y=-0.00013185
MM1212 n33 n113 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.71e-05 $Y=-4.17e-05
MM1181 n6 n97 n113 n6 C5NPMOS w=7.2e-06 l=6e-07 as=1.296e-11 ps=1.8e-05 ad=1.188e-11 pd=1.77e-05 $X=-0.00010335 $Y=-7.68e-05
MM1354 n106 n8 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001437 $Y=5.1e-05
MM1253 n6 n96 n184 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.71e-05 $Y=-4.035e-05
MM1186 n89 n165 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-8.415e-05 $Y=-4.17e-05
MM1326 n6 n108 n146 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001239 $Y=-7.08e-05
MM1361 n163 n64 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001437 $Y=-0.00016245
MM1331 n13 n29 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000129 $Y=2.055e-05
MM1038 n87 n67 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.97e-05 $Y=3.78e-05
MM1185 n178 n86 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-9.135e-05 $Y=-7.68e-05
MM1379 n24 n142 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000159 $Y=2.055e-05
MM1293 n6 n199 n77 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001041 $Y=-4.035e-05
MM1164 n138 n196 n102 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002448 $Y=-5.49e-05
MM1111 n72 n4 n63 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001365 $Y=7.35e-06
MM1180 n6 n165 n11 n6 C5NPMOS w=7.2e-06 l=6e-07 as=1.296e-11 ps=1.8e-05 ad=1.188e-11 pd=1.77e-05 $X=-0.00010335 $Y=-4.53e-05
MM1225 n162 n144 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.935e-05 $Y=-0.00016245
MM1166 n112 n115 n102 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0002499 $Y=-5.49e-05
MM972 n22 n33 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-2.67e-05 $Y=-5.49e-05
MM1406 n158 n138 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002595 $Y=-6.99e-05
MM1098 n71 n146 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000129 $Y=-8.4e-05
MM1165 n125 n7 n48 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00024495 $Y=-3.93e-05
MM1283 n70 n9 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.48e-05 $Y=2.055e-05
MM1256 n82 n114 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.71e-05 $Y=-0.00013185
MM979 n3 n41 n222 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-1.47e-05 $Y=-6.54e-05
MM1153 n7 n75 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00021765 $Y=-3.93e-05
MM1009 n3 n183 n96 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.2e-05 $Y=-5.355e-05
MM1102 n8 n26 n32 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001341 $Y=3.78e-05
MM1147 n112 n84 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000159 $Y=-0.00011445
MM1213 n6 n113 n14 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.71e-05 $Y=-7.68e-05
MM1364 n6 n167 n43 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001488 $Y=-9.15e-06
MM1089 n3 n147 n90 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001239 $Y=-5.355e-05
MM1350 n193 n204 n148 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001365 $Y=-7.08e-05
MM1112 n43 n45 n76 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001365 $Y=-2.235e-05
MM1093 n3 n69 n0 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001239 $Y=-0.00017565
MM1407 n189 n48 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00025965 $Y=-2.61e-05
MM1157 n177 n7 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00022785 $Y=-3.93e-05
MM1059 n30 n190 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001041 $Y=-0.00011445
MM1402 n112 n145 n102 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002499 $Y=-6.99e-05
MM1171 n189 n48 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00025965 $Y=-3.93e-05
MM1128 n3 n167 n43 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001488 $Y=-2.235e-05
MM1388 n196 n75 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002175 $Y=-6.99e-05
MM1084 n56 n164 n107 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001167 $Y=-0.00014505
MM1280 n6 n175 n216 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.97e-05 $Y=-0.00013185
MM1036 n124 n114 n175 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.46e-05 $Y=-0.00014505
MM1187 n86 n165 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-8.415e-05 $Y=-7.68e-05
MM1323 n6 n98 n29 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001239 $Y=2.055e-05
MM1235 n135 n137 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.895e-05 $Y=2.055e-05
MM1076 n132 n105 n107 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001143 $Y=-0.00014505
MM1151 n3 n119 n2 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00021255 $Y=-3.93e-05
MM1373 n212 n95 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001539 $Y=-4.035e-05
MM1264 n175 n114 n12 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.22e-05 $Y=-0.00013185
MM1182 n6 n165 n11 n6 C5NPMOS w=7.2e-06 l=6e-07 as=1.296e-11 ps=1.8e-05 ad=1.188e-11 pd=1.77e-05 $X=-0.00010095 $Y=-4.53e-05
MM1254 n6 n120 n181 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.71e-05 $Y=-7.08e-05
MM1316 n59 n45 n194 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001167 $Y=-9.15e-06
MM1215 n6 n41 n14 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-1.47e-05 $Y=-7.68e-05
MM1335 n126 n18 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000129 $Y=-0.00010125
MM1232 n185 n207 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.175e-05 $Y=-0.00013185
MM1411 n21 n109 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00029925 $Y=-3.735e-05
MM1177 n23 n109 n100 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00030675 $Y=-5.055e-05
MM1386 n145 n119 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002124 $Y=-6.99e-05
MM1206 n5 n54 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-3.63e-05 $Y=-4.17e-05
MM1124 n169 n78 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001437 $Y=-0.00014505
MM1258 n12 n15 n67 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.22e-05 $Y=5.1e-05
MM1041 n3 n50 n154 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.97e-05 $Y=-5.355e-05
MM998 n42 n159 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.895e-05 $Y=3.78e-05
MM1205 n6 n113 n52 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-3.87e-05 $Y=-7.68e-05
MM1163 n182 n177 n48 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00024255 $Y=-3.93e-05
MM1026 n12 n181 n149 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.22e-05 $Y=-8.4e-05
MM1113 n74 n77 n28 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001365 $Y=-5.355e-05
MM1275 n6 n36 n9 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.97e-05 $Y=2.055e-05
MM1039 n9 n36 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.97e-05 $Y=7.35e-06
MM1134 n170 n106 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001539 $Y=3.78e-05
MM1104 n134 n213 n76 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001341 $Y=-2.235e-05
MM1031 n24 n80 n36 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.46e-05 $Y=7.35e-06
MM970 n127 n54 n3 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-3.63e-05 $Y=-5.49e-05
MM1029 n40 n110 n12 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.22e-05 $Y=-0.00017565
MM1413 n100 n21 n23 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00030675 $Y=-3.735e-05
MM1094 n152 n32 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000129 $Y=3.78e-05
MM1327 n6 n208 n18 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001239 $Y=-0.00010125
MM1053 n143 n171 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.48e-05 $Y=-0.00017565
MM1107 n18 n38 n99 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001341 $Y=-0.00011445
MM1241 n6 n162 n139 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.895e-05 $Y=-0.00016245
MM1050 n34 n186 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=9.48e-05 $Y=-8.4e-05
MM1313 n143 n191 n69 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001143 $Y=-0.00016245
MM1384 n6 n168 n124 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000159 $Y=-0.00013185
MM1329 n0 n69 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001239 $Y=-0.00016245
MM1273 n116 n110 n40 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.46e-05 $Y=-0.00016245
MM987 n128 n144 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=1.935e-05 $Y=-0.00011445
MM1062 n3 n121 n26 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001092 $Y=3.78e-05
MM1299 n6 n4 n16 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001092 $Y=2.055e-05
MM1138 n53 n200 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001539 $Y=-8.4e-05
MM984 n218 n144 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=1.935e-05 $Y=-2.235e-05
MM1184 n206 n89 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-9.135e-05 $Y=-4.17e-05
MM1044 n3 n175 n216 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.97e-05 $Y=-0.00014505
MM1207 n6 n41 n52 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-3.63e-05 $Y=-7.68e-05
MM1295 n6 n190 n30 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001041 $Y=-0.00010125
MM1146 n20 n53 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000159 $Y=-8.4e-05
MM1252 n6 n51 n93 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.71e-05 $Y=-9.15e-06
MM1021 n110 n10 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.71e-05 $Y=-0.00017565
MM1148 n124 n168 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000159 $Y=-0.00014505
MM1130 n193 n200 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001488 $Y=-8.4e-05
MM1135 n142 n65 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001539 $Y=7.35e-06
MM1204 n5 n113 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-3.87e-05 $Y=-4.17e-05
MM1028 n175 n82 n12 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.22e-05 $Y=-0.00014505
MM1054 n3 n224 n121 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001041 $Y=3.78e-05
MM1000 n3 n57 n35 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=2.895e-05 $Y=-2.235e-05
MM1086 n32 n174 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001239 $Y=3.78e-05
MM1282 n187 n87 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.48e-05 $Y=5.1e-05
MM1061 n136 n155 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001041 $Y=-0.00017565
MM1173 n23 n189 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00026475 $Y=-3.93e-05
MM1123 n3 n99 n31 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001437 $Y=-0.00011445
MM1376 n6 n169 n168 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001539 $Y=-0.00013185
MM1279 n104 n156 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.97e-05 $Y=-0.00010125
MM994 n103 n62 n201 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=2.175e-05 $Y=-8.4e-05
MM1226 n6 n22 n159 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.175e-05 $Y=5.1e-05
MM1176 n131 n21 n100 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00030435 $Y=-5.055e-05
MM1190 n89 n54 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-7.935e-05 $Y=-4.17e-05
MM1342 n146 n179 n148 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001341 $Y=-7.08e-05
MM1011 n173 n133 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.2e-05 $Y=-0.00011445
MM1234 n42 n159 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.895e-05 $Y=5.1e-05
MM1375 n84 n31 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001539 $Y=-0.00010125
MM954 n217 n54 n3 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-7.935e-05 $Y=-5.49e-05
MM1066 n3 n179 n204 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001092 $Y=-8.4e-05
MM945 n3 n97 n113 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=-0.00010335 $Y=-6.36e-05
MM1010 n3 n55 n120 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=7.2e-05 $Y=-8.4e-05
MM1265 n40 n10 n12 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.22e-05 $Y=-0.00016245
MM1169 n125 n2 n58 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00025245 $Y=-3.93e-05
MM1317 n147 n77 n161 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001167 $Y=-4.035e-05
MM1073 n147 n77 n140 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001143 $Y=-5.355e-05
MM1247 n173 n133 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.2e-05 $Y=-0.00010125
MM1149 n116 n19 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000159 $Y=-0.00017565
MM981 n41 n54 n3 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=-6e-07 $Y=-5.49e-05
MM1314 n174 n121 n152 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001167 $Y=5.1e-05
MM1290 n121 n224 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001041 $Y=5.1e-05
MM1074 n108 n179 n49 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001143 $Y=-8.4e-05
MM1023 n12 n203 n36 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.22e-05 $Y=7.35e-06
MM1288 n172 n216 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.48e-05 $Y=-0.00013185
MM1301 n6 n77 n85 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001092 $Y=-4.035e-05
MM1227 n6 n83 n137 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.175e-05 $Y=2.055e-05
MM993 n94 n206 n215 n3 C5NNMOS w=3.6e-06 l=6e-07 as=2.97e-12 ps=1.05e-05 ad=3.24e-12 pd=1.08e-05 $X=2.175e-05 $Y=-5.355e-05
MM948 n206 n89 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-9.135e-05 $Y=-5.49e-05
MM975 n214 n11 n14 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-1.95e-05 $Y=-6.54e-05
MM1328 n6 n107 n150 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001239 $Y=-0.00013185
MM1366 n193 n200 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001488 $Y=-7.08e-05
MM1217 n6 n54 n41 n6 C5NPMOS w=7.2e-06 l=6e-07 as=1.296e-11 ps=1.8e-05 ad=1.188e-11 pd=1.77e-05 $X=-6e-07 $Y=-4.53e-05
MM1255 n46 n173 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.71e-05 $Y=-0.00010125
MM1139 n3 n31 n84 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001539 $Y=-0.00011445
MM1055 n3 n220 n4 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001041 $Y=7.35e-06
MM1248 n114 n160 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.2e-05 $Y=-0.00013185
MM1140 n168 n169 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001539 $Y=-0.00014505
MM1082 n108 n204 n71 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001167 $Y=-8.4e-05
MM1291 n4 n220 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001041 $Y=2.055e-05
MM1043 n3 n156 n104 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.97e-05 $Y=-0.00011445
MM1239 n133 n39 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.895e-05 $Y=-0.00010125
MM1262 n149 n120 n12 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.22e-05 $Y=-7.08e-05
MM1408 n131 n158 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002646 $Y=-6.99e-05
MM1325 n6 n147 n90 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001239 $Y=-4.035e-05
MM977 n214 n113 n222 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-1.71e-05 $Y=-6.54e-05
MM1222 n103 n144 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.935e-05 $Y=-7.08e-05
MM1276 n211 n27 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=8.97e-05 $Y=-9.15e-06
MM1351 n99 n38 n37 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001365 $Y=-0.00010125
MM1374 n53 n200 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001539 $Y=-7.08e-05
MM1137 n3 n95 n212 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001539 $Y=-5.355e-05
MM1334 n6 n146 n71 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000129 $Y=-7.08e-05
MM1324 n6 n59 n134 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001239 $Y=-9.15e-06
MM1203 n6 n165 n52 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-4.11e-05 $Y=-7.68e-05
MM958 n205 n11 n130 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-6.27e-05 $Y=-5.49e-05
MM1022 n12 n180 n67 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.22e-05 $Y=3.78e-05
MM1297 n136 n155 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001041 $Y=-0.00016245
MM1144 n68 n47 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000159 $Y=-2.235e-05
MM1101 n3 n0 n195 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000129 $Y=-0.00017565
MM1321 n195 n136 n69 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001167 $Y=-0.00016245
MM1395 n24 n118 n182 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00023505 $Y=-2.61e-05
MM1202 n5 n165 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=-4.11e-05 $Y=-4.17e-05
MM1294 n6 n197 n179 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001041 $Y=-7.08e-05
MM1119 n3 n72 n65 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001437 $Y=7.35e-06
MM1236 n6 n57 n35 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.895e-05 $Y=-9.15e-06
MM1228 n6 n17 n57 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=2.175e-05 $Y=-9.15e-06
MM1037 n40 n10 n116 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.46e-05 $Y=-0.00017565
MM1117 n111 n136 n64 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001365 $Y=-0.00017565
MM1345 n0 n136 n64 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001341 $Y=-0.00016245
MM1344 n150 n105 n78 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001341 $Y=-0.00013185
MM1401 n48 n177 n125 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00024495 $Y=-2.61e-05
MM1400 n138 n117 n102 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002448 $Y=-6.99e-05
MM974 n202 n11 n33 n3 C5NNMOS w=5.4e-06 l=6e-07 as=9.72e-12 ps=1.44e-05 ad=8.91e-12 pd=1.41e-05 $X=-1.95e-05 $Y=-5.49e-05
MM1355 n65 n72 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001437 $Y=2.055e-05
MM956 n17 n130 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-6.99e-05 $Y=-5.49e-05
MM1221 n6 n144 n94 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=1.935e-05 $Y=-4.035e-05
MM1287 n73 n104 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=9.48e-05 $Y=-0.00010125
MM1311 n208 n38 n176 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001143 $Y=-0.00010125
MM1302 n6 n179 n204 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001092 $Y=-7.08e-05
MM1242 n15 n42 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.2e-05 $Y=5.1e-05
MM1072 n59 n45 n88 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001143 $Y=-2.235e-05
MM1085 n195 n191 n69 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001167 $Y=-0.00017565
MM1394 n124 n115 n192 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002349 $Y=-6.99e-05
MM1257 n6 n10 n110 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=7.71e-05 $Y=-0.00016245
MM1161 n182 n118 n188 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.00023745 $Y=-3.93e-05
MM1390 n115 n145 n6 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0002226 $Y=-6.99e-05
MM1300 n6 n45 n213 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001092 $Y=-9.15e-06
MM1040 n211 n27 n3 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=8.97e-05 $Y=-2.235e-05
MM1087 n3 n98 n29 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.0001239 $Y=7.35e-06
MM1338 n8 n121 n32 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.0001341 $Y=5.1e-05
MM1414 n6 n100 n25 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.00031185 $Y=-3.735e-05
MM1385 n6 n19 n116 n6 C5NPMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=5.94e-12 pd=1.05e-05 $X=0.000159 $Y=-0.00016245
MM1095 n3 n29 n13 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=0.000129 $Y=7.35e-06
MM957 n3 n129 n207 n3 C5NNMOS w=1.8e-06 l=6e-07 as=2.97e-12 ps=6.9e-06 ad=2.97e-12 pd=6.9e-06 $X=-6.99e-05 $Y=-6.18e-05
.ENDS
