*******************************************************************************
* CDL netlist
*
* Library : buffer_ex
* Top Cell Name: inverter
* View Name: extracted
* Netlist created: 23.Feb.2019 16:18:49
*******************************************************************************

*.SCALE METER
*.GLOBAL VDD VSS

*******************************************************************************
* Library Name: buffer_ex
* Cell Name:    inverter
* View Name:    extracted
*******************************************************************************

.SUBCKT inverter vneg vpos Vin Vout IN
*.PININFO vneg:B vpos:B Vin:B Vout:B IN:B

MM1 vpos Vin Vout vpos C5NPMOS w=1.8e-06 l=6e-07 as=3.78e-12 ps=7.8e-06 ad=3.78e-12 pd=7.8e-06 $X=2.1 $Y=5.4
MM0 vneg Vin Vout vneg C5NNMOS w=1.8e-06 l=6e-07 as=3.78e-12 ps=7.8e-06 ad=3.78e-12 pd=7.8e-06 $X=2.1 $Y=0
.ENDS
