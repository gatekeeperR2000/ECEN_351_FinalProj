*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: inv_8x
* View Name: extracted
* Netlist created: 22.Mar.2019 20:49:56
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    inv_8x
* View Name:    extracted
*******************************************************************************

.SUBCKT inv_8x

MM31 Z A vdd vdd C5NPMOS w=7.2e-06 l=6e-07 as=1.188e-11 ps=1.77e-05 ad=1.296e-11 pd=1.8e-05 $X=11.55 $Y=11.4
MM29 Z A vdd vdd C5NPMOS w=7.2e-06 l=6e-07 as=1.188e-11 ps=1.77e-05 ad=1.296e-11 pd=1.8e-05 $X=6.75 $Y=11.4
MM30 vdd A Z vdd C5NPMOS w=7.2e-06 l=6e-07 as=1.188e-11 ps=1.77e-05 ad=1.296e-11 pd=1.8e-05 $X=9.15 $Y=11.4
MM28 vdd A Z vdd C5NPMOS w=7.2e-06 l=6e-07 as=1.188e-11 ps=1.77e-05 ad=1.296e-11 pd=1.8e-05 $X=4.35 $Y=11.4
MM27 Z A vss vss C5NNMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=6.48e-12 pd=1.08e-05 $X=11.55 $Y=2.4
MM26 vss A Z vss C5NNMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=6.48e-12 pd=1.08e-05 $X=9.15 $Y=2.4
MM25 Z A vss vss C5NNMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=6.48e-12 pd=1.08e-05 $X=6.75 $Y=2.4
MM24 vss A Z vss C5NNMOS w=3.6e-06 l=6e-07 as=5.94e-12 ps=1.05e-05 ad=6.48e-12 pd=1.08e-05 $X=4.35 $Y=2.4
.ENDS
