*******************************************************************************
* CDL netlist
*
* Library : C5N_std_lib
* Top Cell Name: or2_2x
* View Name: schematic
* Netlist created: 23.Mar.2019 20:29:36
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd vss

*******************************************************************************
* Library Name: C5N_std_lib
* Cell Name:    or2_2x
* View Name:    schematic
*******************************************************************************

.SUBCKT or2_2x B A 
*.PININFO Z:O B:I A:I

M4 Z n3 vdd vdd C5NPMOS w=3.6u l=0.6u m=2
M2 n3 B vss vss C5NNMOS w=1.8u l=0.6u m=1
M5 Z n3 vss vss C5NNMOS w=1.8u l=0.6u m=2
M3 n3 B n2 vdd C5NPMOS w=7.2u l=0.6u m=1
M1 n3 A vss vss C5NNMOS w=1.8u l=0.6u m=1
M0 n2 A vdd vdd C5NPMOS w=7.2u l=0.6u m=1
.ENDS

